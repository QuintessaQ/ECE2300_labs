module tffp(RESET, CLK, T);

input RESET; 
input CLK;
input T;

always@(RESET, CLK, T)
begin
	
end